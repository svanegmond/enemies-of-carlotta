From: %(From)s
To: %(To)s
Subject: Prenumeranter på %(list)s
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Här är listan över prenumeranter på listan %(list)s, enligt begäran.

%(addresses)s

Totalt: %(count)s adresser.
