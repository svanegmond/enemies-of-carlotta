From: %(From)s
To: %(To)s
Subject: Adress borttagen från %(list)s
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Hej! 

Det här brevet skickades av epostlistehanteraren som sköter listan

    %(list)s

till listans ägare.

Följande adress har avslutat sin prenumeration på listan:

    %(address)s

Såvida inte något riktigt märkligt pågår är det här brevet bara till
för att informera dig och du behöver inte vidta någon åtgärd.

Tack.