
-- 
Om du vill avsluta prenumerationen, skicka ett brev till
%(local)s-unsubscribe@%(domain)s.
