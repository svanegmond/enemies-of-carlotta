From: %(From)s
To: %(To)s
Subject: Begäran om prenumerantlista för %(list)s nekad
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Tyvärr, du är inte ägaren till listan %(list)s.
