From: %(From)s
To: %(To)s
Subject: Var god vänta på godkännande av prenumerationen på %(list)s
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Hej! 

Det här brevet skickades av epostlistehanteraren som sköter epostlistan
%(list)s.

Du har bekräftat att du vill prenumerera på listan. Prenumerationen är
dock inte öppen för alla, och därför måste listans ägare manuellt 
godkänna din begäran. Det kan ta en stund, så ha tålamod!

För instruktioner om hur man använder epostlistehanteraren, skicka
ett brev till to %(local)s-help@%(domain)s.

Om du har problem, kontakta personerna som äger listan på
%(local)s-owner@%(domain)s.

Tack.
