From: %(From)s
To: %(To)s
Subject: Farväl från %(list)s
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Din prenumeration på %(list)s har härmed avslutats.

För instruktioner om hur man använder epostlistehanteraren, skicka
ett brev till %(local)s-help@%(domain)s.

Om du har problem, kontakta personerna som äger listan på
%(local)s-owner@%(domain)s.

Tack.
