From: %(From)s
To: %(To)s
Subject: Välkommen till %(list)s
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Välkommen till epostlistan %(list)s!

Om du vill avsluta prenumerationen, skicka ett tomt brev till
%(local)s-unsubscribe@%(domain)s.

För instruktioner om hur man använder epostlistehanteraren, skicka
ett brev till %(local)s-help@%(domain)s.

Om du har problem, kontakta personerna som äger listan på
%(local)s-owner@%(domain)s.

Tack.
