From: %(From)s
To: %(To)s
Subject: Prenumerationen på %(list)s avbruten p.g.a. för många studsar
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Hej! 

Du har prenumererat på epostlistan %(list)s.

Tyvärr har post skickad till dig av epostlistehanteraren studsat
så mycket att du har blivit automatiskt borttagen. När problemen
är lösta är du välkommen att prenumerera på nytt.

För instruktioner om hur man använder epostlistehanteraren, skicka
ett brev till to %(local)s-help@%(domain)s.

Om du har problem, kontakta personerna som äger listan på
%(local)s-owner@%(domain)s.

Tack.
