From: %(From)s
To: %(To)s
Subject: Var god vänta på moderering av din postning till %(list)s
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Hej! 

Det här brevet skickades av epostlistehanteraren som sköter epostlistan
%(list)s.

Du, eller någon (kanske en spammer) som föreställer dig, har skickat
ett meddelande till epostlistan. Om det inte var du, var så god och
glöm det här brevet. Om det var du, läs vidare.

Ditt meddelande till listan har skickats till moderatorerna för god-
kännande. Det kan ta ett litet tag. Ha tålamod!

För instruktioner om hur man använder epostlistehanteraren, skicka
ett brev till to %(local)s-help@%(domain)s.

Om du har problem, kontakta personerna som äger listan på
%(local)s-owner@%(domain)s.

Tack.
