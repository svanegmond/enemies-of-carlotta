From: %(From)s
To: %(To)s
Subject: Prenumeration på %(list)s avvisad
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Hej! 

Det här brevet skickades av epostlistehanteraren som sköter epostlistan
%(list)s.

Du försökte prenumerera på listan, men en moderator har avslagit din
begäran. Beklagar.

Om du har problem, kontakta personerna som äger listan på
%(local)s-owner@%(domain)s.

Tack.
