From: %(From)s
To: %(To)s
Subject: Prenumerantlista har ändrats för %(list)s
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Hej! 

Det här brevet skickades av epostlistehanteraren som sköter listan
%(list)s.

För din kännedom: På begäran från en listägare har listan med 
prenumeranter ersatts med en ny.

För instruktioner om hur man använder epostlistehanteraren, skicka
ett brev till to %(local)s-help@%(domain)s.

Om du har problem, kontakta personerna som äger listan på
%(local)s-owner@%(domain)s.

Tack.
