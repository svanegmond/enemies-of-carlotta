From: %(From)s
To: %(To)s
Subject: Du kan inte ställa in prenumerantlistan för %(list)s
Content-type: text/plain; charset=utf-8
MIME-Version: 1.0

Tyvärr, du är inte någon av ägarna till %(list)s.
